`timescale 1ns / 100ps
module top (  /*AUTOARG*/);

  // IOBs

  // PLL

  // Acquisition

  // SDRAM

  // Correlator

  // Output SRAM's

endmodule  // top
